.param W1=10
.param W2=1
