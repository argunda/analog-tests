** sch_path: /home/sai/tt06/analog-tests/inverter/xschem/inverter.sch
**.subckt inverter
XM1 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=W1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=W2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 net1 GND 1.8
V2 IN GND sin(1 1 1e6 0)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/sai/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/sai/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/sai/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/sai/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice




.include guiparams.spice
* These parameters are now set by GUI****
* .param W1=1
* .param W2=1
*****************************************
.control
  reset
  save all
  tran 0.1n 1u
  write inverter.raw
  quit 0
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
